
//module sin(
//input  [10:0]x;
//output [7:0]sinx;
//);
//wire [8:0]x_quatur;
//wire [7:0]tableoutput;

//expand the 1/4 sine to 1/2 sine assume 
//assign x>500?x_quatur = 500-x : x_quatur=x;

//assign sinx = tableoutput;

//if(x[7:0]==255) // if (x == 255)