module  pwm(
		input clk,
		output reg pwm);
		 

	
	
	integer counter;
	integer dut;
	integer div = 5000; // slow down the clock 
	integer r = 0;
	integer delay = 0;
	integer THETA_TMP_COUNTER = 0;
	//integer x;
	
	reg  [9:0] THETA = 10'd0;   // 10 bit, up to 1024
	reg [8:0] THETA_TMP;        //Lower bits of THETA (counting up or counting down)
	reg [9:0] THETA_HLP;        //Helper for reversing lower bits of counting direction for theta
	
	reg [10:0] SINE_TMP;         //Temporary holder for output (two's compliment)
	reg [10:0] SINE_OUT;         //Output Sine in two's compliment
	
always @(posedge clk) begin



    if(r == div ) begin
       THETA = (THETA + 10'b1) % 10'd879; // theta_a is flopped theat 0 to 255  
        r = 1;
		  
		  	//adding delay here 	 
			if(THETA == 10'd0) begin
				THETA_TMP_COUNTER = THETA_TMP_COUNTER + 1;
			end
			else begin
				THETA_TMP_COUNTER = THETA_TMP_COUNTER;
			end

		  //end of delay. 
    end
	 
    else begin
         
		  	if(THETA_TMP_COUNTER == 1) begin
				
			   THETA = 10'd0;
		
				if(delay == 500) begin
					 THETA_TMP_COUNTER = 0;
					 delay = 0;
				end
				else begin 
					delay = delay + 1;
					THETA = 10'd0;
				end 		 
			end	
			else begin
				r = r + 1;	
			end	  
    end
end 
	// pwm generator 
always @(posedge clk) begin
	
	pwm = 1'b1;
	if(counter == 500) begin // Top value, set to setup pwm fre.
		counter = 0;
		pwm = 1'b1; 
	end
	
	else begin
		counter = counter + 1;
		pwm = pwm;
	end
	
	if(counter <= SINE_OUT) // duty cycle value 
		pwm = 1'b1;
	else
		pwm =1'b0;
		
		
end
always @(THETA) begin
	case (THETA)                    			
						
						
		10'd0	:	SINE_TMP	 =	9'd	0	;
		10'd1	:	SINE_TMP	 =	9'd	2	;
		10'd2	:	SINE_TMP	 =	9'd	4	;
		10'd3	:	SINE_TMP	 =	9'd	5	;
		10'd4	:	SINE_TMP	 =	9'd	7	;
		10'd5	:	SINE_TMP	 =	9'd	9	;
		10'd6	:	SINE_TMP	 =	9'd	11	;
		10'd7	:	SINE_TMP	 =	9'd	13	;
		10'd8	:	SINE_TMP	 =	9'd	14	;
		10'd9	:	SINE_TMP	 =	9'd	16	;
		10'd10	:	SINE_TMP	 =	9'd	18	;
		10'd11	:	SINE_TMP	 =	9'd	20	;
		10'd12	:	SINE_TMP	 =	9'd	21	;
		10'd13	:	SINE_TMP	 =	9'd	23	;
		10'd14	:	SINE_TMP	 =	9'd	25	;
		10'd15	:	SINE_TMP	 =	9'd	27	;
		10'd16	:	SINE_TMP	 =	9'd	29	;
		10'd17	:	SINE_TMP	 =	9'd	30	;
		10'd18	:	SINE_TMP	 =	9'd	32	;
		10'd19	:	SINE_TMP	 =	9'd	34	;
		10'd20	:	SINE_TMP	 =	9'd	36	;
		10'd21	:	SINE_TMP	 =	9'd	38	;
		10'd22	:	SINE_TMP	 =	9'd	39	;
		10'd23	:	SINE_TMP	 =	9'd	41	;
		10'd24	:	SINE_TMP	 =	9'd	43	;
		10'd25	:	SINE_TMP	 =	9'd	45	;
		10'd26	:	SINE_TMP	 =	9'd	46	;
		10'd27	:	SINE_TMP	 =	9'd	48	;
		10'd28	:	SINE_TMP	 =	9'd	50	;
		10'd29	:	SINE_TMP	 =	9'd	52	;
		10'd30	:	SINE_TMP	 =	9'd	54	;
		10'd31	:	SINE_TMP	 =	9'd	55	;
		10'd32	:	SINE_TMP	 =	9'd	57	;
		10'd33	:	SINE_TMP	 =	9'd	59	;
		10'd34	:	SINE_TMP	 =	9'd	61	;
		10'd35	:	SINE_TMP	 =	9'd	62	;
		10'd36	:	SINE_TMP	 =	9'd	64	;
		10'd37	:	SINE_TMP	 =	9'd	66	;
		10'd38	:	SINE_TMP	 =	9'd	68	;
		10'd39	:	SINE_TMP	 =	9'd	70	;
		10'd40	:	SINE_TMP	 =	9'd	71	;
		10'd41	:	SINE_TMP	 =	9'd	73	;
		10'd42	:	SINE_TMP	 =	9'd	75	;
		10'd43	:	SINE_TMP	 =	9'd	77	;
		10'd44	:	SINE_TMP	 =	9'd	78	;
		10'd45	:	SINE_TMP	 =	9'd	80	;
		10'd46	:	SINE_TMP	 =	9'd	82	;
		10'd47	:	SINE_TMP	 =	9'd	84	;
		10'd48	:	SINE_TMP	 =	9'd	85	;
		10'd49	:	SINE_TMP	 =	9'd	87	;
		10'd50	:	SINE_TMP	 =	9'd	89	;
		10'd51	:	SINE_TMP	 =	9'd	91	;
		10'd52	:	SINE_TMP	 =	9'd	92	;
		10'd53	:	SINE_TMP	 =	9'd	94	;
		10'd54	:	SINE_TMP	 =	9'd	96	;
		10'd55	:	SINE_TMP	 =	9'd	98	;
		10'd56	:	SINE_TMP	 =	9'd	100	;
		10'd57	:	SINE_TMP	 =	9'd	101	;
		10'd58	:	SINE_TMP	 =	9'd	103	;
		10'd59	:	SINE_TMP	 =	9'd	105	;
		10'd60	:	SINE_TMP	 =	9'd	107	;
		10'd61	:	SINE_TMP	 =	9'd	108	;
		10'd62	:	SINE_TMP	 =	9'd	110	;
		10'd63	:	SINE_TMP	 =	9'd	112	;
		10'd64	:	SINE_TMP	 =	9'd	114	;
		10'd65	:	SINE_TMP	 =	9'd	115	;
		10'd66	:	SINE_TMP	 =	9'd	117	;
		10'd67	:	SINE_TMP	 =	9'd	119	;
		10'd68	:	SINE_TMP	 =	9'd	120	;
		10'd69	:	SINE_TMP	 =	9'd	122	;
		10'd70	:	SINE_TMP	 =	9'd	124	;
		10'd71	:	SINE_TMP	 =	9'd	126	;
		10'd72	:	SINE_TMP	 =	9'd	127	;
		10'd73	:	SINE_TMP	 =	9'd	129	;
		10'd74	:	SINE_TMP	 =	9'd	131	;
		10'd75	:	SINE_TMP	 =	9'd	133	;
		10'd76	:	SINE_TMP	 =	9'd	134	;
		10'd77	:	SINE_TMP	 =	9'd	136	;
		10'd78	:	SINE_TMP	 =	9'd	138	;
		10'd79	:	SINE_TMP	 =	9'd	139	;
		10'd80	:	SINE_TMP	 =	9'd	141	;
		10'd81	:	SINE_TMP	 =	9'd	143	;
		10'd82	:	SINE_TMP	 =	9'd	145	;
		10'd83	:	SINE_TMP	 =	9'd	146	;
		10'd84	:	SINE_TMP	 =	9'd	148	;
		10'd85	:	SINE_TMP	 =	9'd	150	;
		10'd86	:	SINE_TMP	 =	9'd	151	;
		10'd87	:	SINE_TMP	 =	9'd	153	;
		10'd88	:	SINE_TMP	 =	9'd	155	;
		10'd89	:	SINE_TMP	 =	9'd	157	;
		10'd90	:	SINE_TMP	 =	9'd	158	;
		10'd91	:	SINE_TMP	 =	9'd	160	;
		10'd92	:	SINE_TMP	 =	9'd	162	;
		10'd93	:	SINE_TMP	 =	9'd	163	;
		10'd94	:	SINE_TMP	 =	9'd	165	;
		10'd95	:	SINE_TMP	 =	9'd	167	;
		10'd96	:	SINE_TMP	 =	9'd	168	;
		10'd97	:	SINE_TMP	 =	9'd	170	;
		10'd98	:	SINE_TMP	 =	9'd	172	;
		10'd99	:	SINE_TMP	 =	9'd	173	;
		10'd100	:	SINE_TMP	 =	9'd	175	;
		10'd101	:	SINE_TMP	 =	9'd	177	;
		10'd102	:	SINE_TMP	 =	9'd	178	;
		10'd103	:	SINE_TMP	 =	9'd	180	;
		10'd104	:	SINE_TMP	 =	9'd	182	;
		10'd105	:	SINE_TMP	 =	9'd	183	;
		10'd106	:	SINE_TMP	 =	9'd	185	;
		10'd107	:	SINE_TMP	 =	9'd	187	;
		10'd108	:	SINE_TMP	 =	9'd	188	;
		10'd109	:	SINE_TMP	 =	9'd	190	;
		10'd110	:	SINE_TMP	 =	9'd	192	;
		10'd111	:	SINE_TMP	 =	9'd	193	;
		10'd112	:	SINE_TMP	 =	9'd	195	;
		10'd113	:	SINE_TMP	 =	9'd	197	;
		10'd114	:	SINE_TMP	 =	9'd	198	;
		10'd115	:	SINE_TMP	 =	9'd	200	;
		10'd116	:	SINE_TMP	 =	9'd	202	;
		10'd117	:	SINE_TMP	 =	9'd	203	;
		10'd118	:	SINE_TMP	 =	9'd	205	;
		10'd119	:	SINE_TMP	 =	9'd	207	;
		10'd120	:	SINE_TMP	 =	9'd	208	;
		10'd121	:	SINE_TMP	 =	9'd	210	;
		10'd122	:	SINE_TMP	 =	9'd	211	;
		10'd123	:	SINE_TMP	 =	9'd	213	;
		10'd124	:	SINE_TMP	 =	9'd	215	;
		10'd125	:	SINE_TMP	 =	9'd	216	;
		10'd126	:	SINE_TMP	 =	9'd	218	;
		10'd127	:	SINE_TMP	 =	9'd	219	;
		10'd128	:	SINE_TMP	 =	9'd	221	;
		10'd129	:	SINE_TMP	 =	9'd	223	;
		10'd130	:	SINE_TMP	 =	9'd	224	;
		10'd131	:	SINE_TMP	 =	9'd	226	;
		10'd132	:	SINE_TMP	 =	9'd	227	;
		10'd133	:	SINE_TMP	 =	9'd	229	;
		10'd134	:	SINE_TMP	 =	9'd	231	;
		10'd135	:	SINE_TMP	 =	9'd	232	;
		10'd136	:	SINE_TMP	 =	9'd	234	;
		10'd137	:	SINE_TMP	 =	9'd	235	;
		10'd138	:	SINE_TMP	 =	9'd	237	;
		10'd139	:	SINE_TMP	 =	9'd	239	;
		10'd140	:	SINE_TMP	 =	9'd	240	;
		10'd141	:	SINE_TMP	 =	9'd	242	;
		10'd142	:	SINE_TMP	 =	9'd	243	;
		10'd143	:	SINE_TMP	 =	9'd	245	;
		10'd144	:	SINE_TMP	 =	9'd	246	;
		10'd145	:	SINE_TMP	 =	9'd	248	;
		10'd146	:	SINE_TMP	 =	9'd	249	;
		10'd147	:	SINE_TMP	 =	9'd	251	;
		10'd148	:	SINE_TMP	 =	9'd	253	;
		10'd149	:	SINE_TMP	 =	9'd	254	;
		10'd150	:	SINE_TMP	 =	9'd	256	;
		10'd151	:	SINE_TMP	 =	9'd	257	;
		10'd152	:	SINE_TMP	 =	9'd	259	;
		10'd153	:	SINE_TMP	 =	9'd	260	;
		10'd154	:	SINE_TMP	 =	9'd	262	;
		10'd155	:	SINE_TMP	 =	9'd	263	;
		10'd156	:	SINE_TMP	 =	9'd	265	;
		10'd157	:	SINE_TMP	 =	9'd	266	;
		10'd158	:	SINE_TMP	 =	9'd	268	;
		10'd159	:	SINE_TMP	 =	9'd	269	;
		10'd160	:	SINE_TMP	 =	9'd	271	;
		10'd161	:	SINE_TMP	 =	9'd	272	;
		10'd162	:	SINE_TMP	 =	9'd	274	;
		10'd163	:	SINE_TMP	 =	9'd	275	;
		10'd164	:	SINE_TMP	 =	9'd	277	;
		10'd165	:	SINE_TMP	 =	9'd	278	;
		10'd166	:	SINE_TMP	 =	9'd	280	;
		10'd167	:	SINE_TMP	 =	9'd	281	;
		10'd168	:	SINE_TMP	 =	9'd	283	;
		10'd169	:	SINE_TMP	 =	9'd	284	;
		10'd170	:	SINE_TMP	 =	9'd	286	;
		10'd171	:	SINE_TMP	 =	9'd	287	;
		10'd172	:	SINE_TMP	 =	9'd	289	;
		10'd173	:	SINE_TMP	 =	9'd	290	;
		10'd174	:	SINE_TMP	 =	9'd	292	;
		10'd175	:	SINE_TMP	 =	9'd	293	;
		10'd176	:	SINE_TMP	 =	9'd	294	;
		10'd177	:	SINE_TMP	 =	9'd	296	;
		10'd178	:	SINE_TMP	 =	9'd	297	;
		10'd179	:	SINE_TMP	 =	9'd	299	;
		10'd180	:	SINE_TMP	 =	9'd	300	;
		10'd181	:	SINE_TMP	 =	9'd	302	;
		10'd182	:	SINE_TMP	 =	9'd	303	;
		10'd183	:	SINE_TMP	 =	9'd	304	;
		10'd184	:	SINE_TMP	 =	9'd	306	;
		10'd185	:	SINE_TMP	 =	9'd	307	;
		10'd186	:	SINE_TMP	 =	9'd	309	;
		10'd187	:	SINE_TMP	 =	9'd	310	;
		10'd188	:	SINE_TMP	 =	9'd	312	;
		10'd189	:	SINE_TMP	 =	9'd	313	;
		10'd190	:	SINE_TMP	 =	9'd	314	;
		10'd191	:	SINE_TMP	 =	9'd	316	;
		10'd192	:	SINE_TMP	 =	9'd	317	;
		10'd193	:	SINE_TMP	 =	9'd	318	;
		10'd194	:	SINE_TMP	 =	9'd	320	;
		10'd195	:	SINE_TMP	 =	9'd	321	;
		10'd196	:	SINE_TMP	 =	9'd	323	;
		10'd197	:	SINE_TMP	 =	9'd	324	;
		10'd198	:	SINE_TMP	 =	9'd	325	;
		10'd199	:	SINE_TMP	 =	9'd	327	;
		10'd200	:	SINE_TMP	 =	9'd	328	;
		10'd201	:	SINE_TMP	 =	9'd	329	;
		10'd202	:	SINE_TMP	 =	9'd	331	;
		10'd203	:	SINE_TMP	 =	9'd	332	;
		10'd204	:	SINE_TMP	 =	9'd	333	;
		10'd205	:	SINE_TMP	 =	9'd	335	;
		10'd206	:	SINE_TMP	 =	9'd	336	;
		10'd207	:	SINE_TMP	 =	9'd	337	;
		10'd208	:	SINE_TMP	 =	9'd	339	;
		10'd209	:	SINE_TMP	 =	9'd	340	;
		10'd210	:	SINE_TMP	 =	9'd	341	;
		10'd211	:	SINE_TMP	 =	9'd	343	;
		10'd212	:	SINE_TMP	 =	9'd	344	;
		10'd213	:	SINE_TMP	 =	9'd	345	;
		10'd214	:	SINE_TMP	 =	9'd	347	;
		10'd215	:	SINE_TMP	 =	9'd	348	;
		10'd216	:	SINE_TMP	 =	9'd	349	;
		10'd217	:	SINE_TMP	 =	9'd	350	;
		10'd218	:	SINE_TMP	 =	9'd	352	;
		10'd219	:	SINE_TMP	 =	9'd	353	;
		10'd220	:	SINE_TMP	 =	9'd	354	;
		10'd221	:	SINE_TMP	 =	9'd	355	;
		10'd222	:	SINE_TMP	 =	9'd	357	;
		10'd223	:	SINE_TMP	 =	9'd	358	;
		10'd224	:	SINE_TMP	 =	9'd	359	;
		10'd225	:	SINE_TMP	 =	9'd	360	;
		10'd226	:	SINE_TMP	 =	9'd	362	;
		10'd227	:	SINE_TMP	 =	9'd	363	;
		10'd228	:	SINE_TMP	 =	9'd	364	;
		10'd229	:	SINE_TMP	 =	9'd	365	;
		10'd230	:	SINE_TMP	 =	9'd	367	;
		10'd231	:	SINE_TMP	 =	9'd	368	;
		10'd232	:	SINE_TMP	 =	9'd	369	;
		10'd233	:	SINE_TMP	 =	9'd	370	;
		10'd234	:	SINE_TMP	 =	9'd	371	;
		10'd235	:	SINE_TMP	 =	9'd	373	;
		10'd236	:	SINE_TMP	 =	9'd	374	;
		10'd237	:	SINE_TMP	 =	9'd	375	;
		10'd238	:	SINE_TMP	 =	9'd	376	;
		10'd239	:	SINE_TMP	 =	9'd	377	;
		10'd240	:	SINE_TMP	 =	9'd	379	;
		10'd241	:	SINE_TMP	 =	9'd	380	;
		10'd242	:	SINE_TMP	 =	9'd	381	;
		10'd243	:	SINE_TMP	 =	9'd	382	;
		10'd244	:	SINE_TMP	 =	9'd	383	;
		10'd245	:	SINE_TMP	 =	9'd	384	;
		10'd246	:	SINE_TMP	 =	9'd	385	;
		10'd247	:	SINE_TMP	 =	9'd	387	;
		10'd248	:	SINE_TMP	 =	9'd	388	;
		10'd249	:	SINE_TMP	 =	9'd	389	;
		10'd250	:	SINE_TMP	 =	9'd	390	;
		10'd251	:	SINE_TMP	 =	9'd	391	;
		10'd252	:	SINE_TMP	 =	9'd	392	;
		10'd253	:	SINE_TMP	 =	9'd	393	;
		10'd254	:	SINE_TMP	 =	9'd	394	;
		10'd255	:	SINE_TMP	 =	9'd	395	;
		10'd256	:	SINE_TMP	 =	9'd	397	;
		10'd257	:	SINE_TMP	 =	9'd	398	;
		10'd258	:	SINE_TMP	 =	9'd	399	;
		10'd259	:	SINE_TMP	 =	9'd	400	;
		10'd260	:	SINE_TMP	 =	9'd	401	;
		10'd261	:	SINE_TMP	 =	9'd	402	;
		10'd262	:	SINE_TMP	 =	9'd	403	;
		10'd263	:	SINE_TMP	 =	9'd	404	;
		10'd264	:	SINE_TMP	 =	9'd	405	;
		10'd265	:	SINE_TMP	 =	9'd	406	;
		10'd266	:	SINE_TMP	 =	9'd	407	;
		10'd267	:	SINE_TMP	 =	9'd	408	;
		10'd268	:	SINE_TMP	 =	9'd	409	;
		10'd269	:	SINE_TMP	 =	9'd	410	;
		10'd270	:	SINE_TMP	 =	9'd	411	;
		10'd271	:	SINE_TMP	 =	9'd	412	;
		10'd272	:	SINE_TMP	 =	9'd	413	;
		10'd273	:	SINE_TMP	 =	9'd	414	;
		10'd274	:	SINE_TMP	 =	9'd	415	;
		10'd275	:	SINE_TMP	 =	9'd	416	;
		10'd276	:	SINE_TMP	 =	9'd	417	;
		10'd277	:	SINE_TMP	 =	9'd	418	;
		10'd278	:	SINE_TMP	 =	9'd	419	;
		10'd279	:	SINE_TMP	 =	9'd	420	;
		10'd280	:	SINE_TMP	 =	9'd	421	;
		10'd281	:	SINE_TMP	 =	9'd	422	;
		10'd282	:	SINE_TMP	 =	9'd	423	;
		10'd283	:	SINE_TMP	 =	9'd	424	;
		10'd284	:	SINE_TMP	 =	9'd	425	;
		10'd285	:	SINE_TMP	 =	9'd	426	;
		10'd286	:	SINE_TMP	 =	9'd	427	;
		10'd287	:	SINE_TMP	 =	9'd	428	;
		10'd288	:	SINE_TMP	 =	9'd	429	;
		10'd289	:	SINE_TMP	 =	9'd	430	;
		10'd290	:	SINE_TMP	 =	9'd	431	;
		10'd291	:	SINE_TMP	 =	9'd	432	;
		10'd292	:	SINE_TMP	 =	9'd	432	;
		10'd293	:	SINE_TMP	 =	9'd	433	;
		10'd294	:	SINE_TMP	 =	9'd	434	;
		10'd295	:	SINE_TMP	 =	9'd	435	;
		10'd296	:	SINE_TMP	 =	9'd	436	;
		10'd297	:	SINE_TMP	 =	9'd	437	;
		10'd298	:	SINE_TMP	 =	9'd	438	;
		10'd299	:	SINE_TMP	 =	9'd	439	;
		10'd300	:	SINE_TMP	 =	9'd	439	;
		10'd301	:	SINE_TMP	 =	9'd	440	;
		10'd302	:	SINE_TMP	 =	9'd	441	;
		10'd303	:	SINE_TMP	 =	9'd	442	;
		10'd304	:	SINE_TMP	 =	9'd	443	;
		10'd305	:	SINE_TMP	 =	9'd	444	;
		10'd306	:	SINE_TMP	 =	9'd	444	;
		10'd307	:	SINE_TMP	 =	9'd	445	;
		10'd308	:	SINE_TMP	 =	9'd	446	;
		10'd309	:	SINE_TMP	 =	9'd	447	;
		10'd310	:	SINE_TMP	 =	9'd	448	;
		10'd311	:	SINE_TMP	 =	9'd	448	;
		10'd312	:	SINE_TMP	 =	9'd	449	;
		10'd313	:	SINE_TMP	 =	9'd	450	;
		10'd314	:	SINE_TMP	 =	9'd	451	;
		10'd315	:	SINE_TMP	 =	9'd	452	;
		10'd316	:	SINE_TMP	 =	9'd	452	;
		10'd317	:	SINE_TMP	 =	9'd	453	;
		10'd318	:	SINE_TMP	 =	9'd	454	;
		10'd319	:	SINE_TMP	 =	9'd	455	;
		10'd320	:	SINE_TMP	 =	9'd	455	;
		10'd321	:	SINE_TMP	 =	9'd	456	;
		10'd322	:	SINE_TMP	 =	9'd	457	;
		10'd323	:	SINE_TMP	 =	9'd	458	;
		10'd324	:	SINE_TMP	 =	9'd	458	;
		10'd325	:	SINE_TMP	 =	9'd	459	;
		10'd326	:	SINE_TMP	 =	9'd	460	;
		10'd327	:	SINE_TMP	 =	9'd	460	;
		10'd328	:	SINE_TMP	 =	9'd	461	;
		10'd329	:	SINE_TMP	 =	9'd	462	;
		10'd330	:	SINE_TMP	 =	9'd	462	;
		10'd331	:	SINE_TMP	 =	9'd	463	;
		10'd332	:	SINE_TMP	 =	9'd	464	;
		10'd333	:	SINE_TMP	 =	9'd	464	;
		10'd334	:	SINE_TMP	 =	9'd	465	;
		10'd335	:	SINE_TMP	 =	9'd	466	;
		10'd336	:	SINE_TMP	 =	9'd	466	;
		10'd337	:	SINE_TMP	 =	9'd	467	;
		10'd338	:	SINE_TMP	 =	9'd	468	;
		10'd339	:	SINE_TMP	 =	9'd	468	;
		10'd340	:	SINE_TMP	 =	9'd	469	;
		10'd341	:	SINE_TMP	 =	9'd	470	;
		10'd342	:	SINE_TMP	 =	9'd	470	;
		10'd343	:	SINE_TMP	 =	9'd	471	;
		10'd344	:	SINE_TMP	 =	9'd	471	;
		10'd345	:	SINE_TMP	 =	9'd	472	;
		10'd346	:	SINE_TMP	 =	9'd	473	;
		10'd347	:	SINE_TMP	 =	9'd	473	;
		10'd348	:	SINE_TMP	 =	9'd	474	;
		10'd349	:	SINE_TMP	 =	9'd	474	;
		10'd350	:	SINE_TMP	 =	9'd	475	;
		10'd351	:	SINE_TMP	 =	9'd	475	;
		10'd352	:	SINE_TMP	 =	9'd	476	;
		10'd353	:	SINE_TMP	 =	9'd	477	;
		10'd354	:	SINE_TMP	 =	9'd	477	;
		10'd355	:	SINE_TMP	 =	9'd	478	;
		10'd356	:	SINE_TMP	 =	9'd	478	;
		10'd357	:	SINE_TMP	 =	9'd	479	;
		10'd358	:	SINE_TMP	 =	9'd	479	;
		10'd359	:	SINE_TMP	 =	9'd	480	;
		10'd360	:	SINE_TMP	 =	9'd	480	;
		10'd361	:	SINE_TMP	 =	9'd	481	;
		10'd362	:	SINE_TMP	 =	9'd	481	;
		10'd363	:	SINE_TMP	 =	9'd	482	;
		10'd364	:	SINE_TMP	 =	9'd	482	;
		10'd365	:	SINE_TMP	 =	9'd	483	;
		10'd366	:	SINE_TMP	 =	9'd	483	;
		10'd367	:	SINE_TMP	 =	9'd	483	;
		10'd368	:	SINE_TMP	 =	9'd	484	;
		10'd369	:	SINE_TMP	 =	9'd	484	;
		10'd370	:	SINE_TMP	 =	9'd	485	;
		10'd371	:	SINE_TMP	 =	9'd	485	;
		10'd372	:	SINE_TMP	 =	9'd	486	;
		10'd373	:	SINE_TMP	 =	9'd	486	;
		10'd374	:	SINE_TMP	 =	9'd	487	;
		10'd375	:	SINE_TMP	 =	9'd	487	;
		10'd376	:	SINE_TMP	 =	9'd	487	;
		10'd377	:	SINE_TMP	 =	9'd	488	;
		10'd378	:	SINE_TMP	 =	9'd	488	;
		10'd379	:	SINE_TMP	 =	9'd	489	;
		10'd380	:	SINE_TMP	 =	9'd	489	;
		10'd381	:	SINE_TMP	 =	9'd	489	;
		10'd382	:	SINE_TMP	 =	9'd	490	;
		10'd383	:	SINE_TMP	 =	9'd	490	;
		10'd384	:	SINE_TMP	 =	9'd	490	;
		10'd385	:	SINE_TMP	 =	9'd	491	;
		10'd386	:	SINE_TMP	 =	9'd	491	;
		10'd387	:	SINE_TMP	 =	9'd	491	;
		10'd388	:	SINE_TMP	 =	9'd	492	;
		10'd389	:	SINE_TMP	 =	9'd	492	;
		10'd390	:	SINE_TMP	 =	9'd	492	;
		10'd391	:	SINE_TMP	 =	9'd	493	;
		10'd392	:	SINE_TMP	 =	9'd	493	;
		10'd393	:	SINE_TMP	 =	9'd	493	;
		10'd394	:	SINE_TMP	 =	9'd	494	;
		10'd395	:	SINE_TMP	 =	9'd	494	;
		10'd396	:	SINE_TMP	 =	9'd	494	;
		10'd397	:	SINE_TMP	 =	9'd	494	;
		10'd398	:	SINE_TMP	 =	9'd	495	;
		10'd399	:	SINE_TMP	 =	9'd	495	;
		10'd400	:	SINE_TMP	 =	9'd	495	;
		10'd401	:	SINE_TMP	 =	9'd	495	;
		10'd402	:	SINE_TMP	 =	9'd	496	;
		10'd403	:	SINE_TMP	 =	9'd	496	;
		10'd404	:	SINE_TMP	 =	9'd	496	;
		10'd405	:	SINE_TMP	 =	9'd	496	;
		10'd406	:	SINE_TMP	 =	9'd	497	;
		10'd407	:	SINE_TMP	 =	9'd	497	;
		10'd408	:	SINE_TMP	 =	9'd	497	;
		10'd409	:	SINE_TMP	 =	9'd	497	;
		10'd410	:	SINE_TMP	 =	9'd	497	;
		10'd411	:	SINE_TMP	 =	9'd	497	;
		10'd412	:	SINE_TMP	 =	9'd	498	;
		10'd413	:	SINE_TMP	 =	9'd	498	;
		10'd414	:	SINE_TMP	 =	9'd	498	;
		10'd415	:	SINE_TMP	 =	9'd	498	;
		10'd416	:	SINE_TMP	 =	9'd	498	;
		10'd417	:	SINE_TMP	 =	9'd	498	;
		10'd418	:	SINE_TMP	 =	9'd	499	;
		10'd419	:	SINE_TMP	 =	9'd	499	;
		10'd420	:	SINE_TMP	 =	9'd	499	;
		10'd421	:	SINE_TMP	 =	9'd	499	;
		10'd422	:	SINE_TMP	 =	9'd	499	;
		10'd423	:	SINE_TMP	 =	9'd	499	;
		10'd424	:	SINE_TMP	 =	9'd	499	;
		10'd425	:	SINE_TMP	 =	9'd	499	;
		10'd426	:	SINE_TMP	 =	9'd	499	;
		10'd427	:	SINE_TMP	 =	9'd	500	;
		10'd428	:	SINE_TMP	 =	9'd	500	;
		10'd429	:	SINE_TMP	 =	9'd	500	;
		10'd430	:	SINE_TMP	 =	9'd	500	;
		10'd431	:	SINE_TMP	 =	9'd	500	;
		10'd432	:	SINE_TMP	 =	9'd	500	;
		10'd433	:	SINE_TMP	 =	9'd	500	;
		10'd434	:	SINE_TMP	 =	9'd	500	;
		10'd435	:	SINE_TMP	 =	9'd	500	;
		10'd436	:	SINE_TMP	 =	9'd	500	;
		10'd437	:	SINE_TMP	 =	9'd	500	;
		10'd438	:	SINE_TMP	 =	9'd	500	;
		10'd439	:	SINE_TMP	 =	9'd	500	;
		10'd440	:	SINE_TMP	 =	9'd	500	;
		10'd441	:	SINE_TMP	 =	9'd	500	;
		10'd442	:	SINE_TMP	 =	9'd	500	;
		10'd443	:	SINE_TMP	 =	9'd	500	;
		10'd444	:	SINE_TMP	 =	9'd	500	;
		10'd445	:	SINE_TMP	 =	9'd	500	;
		10'd446	:	SINE_TMP	 =	9'd	500	;
		10'd447	:	SINE_TMP	 =	9'd	500	;
		10'd448	:	SINE_TMP	 =	9'd	500	;
		10'd449	:	SINE_TMP	 =	9'd	500	;
		10'd450	:	SINE_TMP	 =	9'd	500	;
		10'd451	:	SINE_TMP	 =	9'd	500	;
		10'd452	:	SINE_TMP	 =	9'd	499	;
		10'd453	:	SINE_TMP	 =	9'd	499	;
		10'd454	:	SINE_TMP	 =	9'd	499	;
		10'd455	:	SINE_TMP	 =	9'd	499	;
		10'd456	:	SINE_TMP	 =	9'd	499	;
		10'd457	:	SINE_TMP	 =	9'd	499	;
		10'd458	:	SINE_TMP	 =	9'd	499	;
		10'd459	:	SINE_TMP	 =	9'd	499	;
		10'd460	:	SINE_TMP	 =	9'd	499	;
		10'd461	:	SINE_TMP	 =	9'd	498	;
		10'd462	:	SINE_TMP	 =	9'd	498	;
		10'd463	:	SINE_TMP	 =	9'd	498	;
		10'd464	:	SINE_TMP	 =	9'd	498	;
		10'd465	:	SINE_TMP	 =	9'd	498	;
		10'd466	:	SINE_TMP	 =	9'd	498	;
		10'd467	:	SINE_TMP	 =	9'd	497	;
		10'd468	:	SINE_TMP	 =	9'd	497	;
		10'd469	:	SINE_TMP	 =	9'd	497	;
		10'd470	:	SINE_TMP	 =	9'd	497	;
		10'd471	:	SINE_TMP	 =	9'd	497	;
		10'd472	:	SINE_TMP	 =	9'd	497	;
		10'd473	:	SINE_TMP	 =	9'd	496	;
		10'd474	:	SINE_TMP	 =	9'd	496	;
		10'd475	:	SINE_TMP	 =	9'd	496	;
		10'd476	:	SINE_TMP	 =	9'd	496	;
		10'd477	:	SINE_TMP	 =	9'd	495	;
		10'd478	:	SINE_TMP	 =	9'd	495	;
		10'd479	:	SINE_TMP	 =	9'd	495	;
		10'd480	:	SINE_TMP	 =	9'd	495	;
		10'd481	:	SINE_TMP	 =	9'd	494	;
		10'd482	:	SINE_TMP	 =	9'd	494	;
		10'd483	:	SINE_TMP	 =	9'd	494	;
		10'd484	:	SINE_TMP	 =	9'd	494	;
		10'd485	:	SINE_TMP	 =	9'd	493	;
		10'd486	:	SINE_TMP	 =	9'd	493	;
		10'd487	:	SINE_TMP	 =	9'd	493	;
		10'd488	:	SINE_TMP	 =	9'd	492	;
		10'd489	:	SINE_TMP	 =	9'd	492	;
		10'd490	:	SINE_TMP	 =	9'd	492	;
		10'd491	:	SINE_TMP	 =	9'd	491	;
		10'd492	:	SINE_TMP	 =	9'd	491	;
		10'd493	:	SINE_TMP	 =	9'd	491	;
		10'd494	:	SINE_TMP	 =	9'd	490	;
		10'd495	:	SINE_TMP	 =	9'd	490	;
		10'd496	:	SINE_TMP	 =	9'd	490	;
		10'd497	:	SINE_TMP	 =	9'd	489	;
		10'd498	:	SINE_TMP	 =	9'd	489	;
		10'd499	:	SINE_TMP	 =	9'd	489	;
		10'd500	:	SINE_TMP	 =	9'd	488	;
		10'd501	:	SINE_TMP	 =	9'd	488	;
		10'd502	:	SINE_TMP	 =	9'd	487	;
		10'd503	:	SINE_TMP	 =	9'd	487	;
		10'd504	:	SINE_TMP	 =	9'd	487	;
		10'd505	:	SINE_TMP	 =	9'd	486	;
		10'd506	:	SINE_TMP	 =	9'd	486	;
		10'd507	:	SINE_TMP	 =	9'd	485	;
		10'd508	:	SINE_TMP	 =	9'd	485	;
		10'd509	:	SINE_TMP	 =	9'd	484	;
		10'd510	:	SINE_TMP	 =	9'd	484	;
		10'd511	:	SINE_TMP	 =	9'd	483	;
		10'd512	:	SINE_TMP	 =	9'd	483	;
		10'd513	:	SINE_TMP	 =	9'd	483	;
		10'd514	:	SINE_TMP	 =	9'd	482	;
		10'd515	:	SINE_TMP	 =	9'd	482	;
		10'd516	:	SINE_TMP	 =	9'd	481	;
		10'd517	:	SINE_TMP	 =	9'd	481	;
		10'd518	:	SINE_TMP	 =	9'd	480	;
		10'd519	:	SINE_TMP	 =	9'd	480	;
		10'd520	:	SINE_TMP	 =	9'd	479	;
		10'd521	:	SINE_TMP	 =	9'd	479	;
		10'd522	:	SINE_TMP	 =	9'd	478	;
		10'd523	:	SINE_TMP	 =	9'd	478	;
		10'd524	:	SINE_TMP	 =	9'd	477	;
		10'd525	:	SINE_TMP	 =	9'd	477	;
		10'd526	:	SINE_TMP	 =	9'd	476	;
		10'd527	:	SINE_TMP	 =	9'd	475	;
		10'd528	:	SINE_TMP	 =	9'd	475	;
		10'd529	:	SINE_TMP	 =	9'd	474	;
		10'd530	:	SINE_TMP	 =	9'd	474	;
		10'd531	:	SINE_TMP	 =	9'd	473	;
		10'd532	:	SINE_TMP	 =	9'd	473	;
		10'd533	:	SINE_TMP	 =	9'd	472	;
		10'd534	:	SINE_TMP	 =	9'd	471	;
		10'd535	:	SINE_TMP	 =	9'd	471	;
		10'd536	:	SINE_TMP	 =	9'd	470	;
		10'd537	:	SINE_TMP	 =	9'd	470	;
		10'd538	:	SINE_TMP	 =	9'd	469	;
		10'd539	:	SINE_TMP	 =	9'd	468	;
		10'd540	:	SINE_TMP	 =	9'd	468	;
		10'd541	:	SINE_TMP	 =	9'd	467	;
		10'd542	:	SINE_TMP	 =	9'd	466	;
		10'd543	:	SINE_TMP	 =	9'd	466	;
		10'd544	:	SINE_TMP	 =	9'd	465	;
		10'd545	:	SINE_TMP	 =	9'd	464	;
		10'd546	:	SINE_TMP	 =	9'd	464	;
		10'd547	:	SINE_TMP	 =	9'd	463	;
		10'd548	:	SINE_TMP	 =	9'd	462	;
		10'd549	:	SINE_TMP	 =	9'd	462	;
		10'd550	:	SINE_TMP	 =	9'd	461	;
		10'd551	:	SINE_TMP	 =	9'd	460	;
		10'd552	:	SINE_TMP	 =	9'd	460	;
		10'd553	:	SINE_TMP	 =	9'd	459	;
		10'd554	:	SINE_TMP	 =	9'd	458	;
		10'd555	:	SINE_TMP	 =	9'd	458	;
		10'd556	:	SINE_TMP	 =	9'd	457	;
		10'd557	:	SINE_TMP	 =	9'd	456	;
		10'd558	:	SINE_TMP	 =	9'd	455	;
		10'd559	:	SINE_TMP	 =	9'd	455	;
		10'd560	:	SINE_TMP	 =	9'd	454	;
		10'd561	:	SINE_TMP	 =	9'd	453	;
		10'd562	:	SINE_TMP	 =	9'd	452	;
		10'd563	:	SINE_TMP	 =	9'd	452	;
		10'd564	:	SINE_TMP	 =	9'd	451	;
		10'd565	:	SINE_TMP	 =	9'd	450	;
		10'd566	:	SINE_TMP	 =	9'd	449	;
		10'd567	:	SINE_TMP	 =	9'd	448	;
		10'd568	:	SINE_TMP	 =	9'd	448	;
		10'd569	:	SINE_TMP	 =	9'd	447	;
		10'd570	:	SINE_TMP	 =	9'd	446	;
		10'd571	:	SINE_TMP	 =	9'd	445	;
		10'd572	:	SINE_TMP	 =	9'd	444	;
		10'd573	:	SINE_TMP	 =	9'd	444	;
		10'd574	:	SINE_TMP	 =	9'd	443	;
		10'd575	:	SINE_TMP	 =	9'd	442	;
		10'd576	:	SINE_TMP	 =	9'd	441	;
		10'd577	:	SINE_TMP	 =	9'd	440	;
		10'd578	:	SINE_TMP	 =	9'd	439	;
		10'd579	:	SINE_TMP	 =	9'd	439	;
		10'd580	:	SINE_TMP	 =	9'd	438	;
		10'd581	:	SINE_TMP	 =	9'd	437	;
		10'd582	:	SINE_TMP	 =	9'd	436	;
		10'd583	:	SINE_TMP	 =	9'd	435	;
		10'd584	:	SINE_TMP	 =	9'd	434	;
		10'd585	:	SINE_TMP	 =	9'd	433	;
		10'd586	:	SINE_TMP	 =	9'd	432	;
		10'd587	:	SINE_TMP	 =	9'd	432	;
		10'd588	:	SINE_TMP	 =	9'd	431	;
		10'd589	:	SINE_TMP	 =	9'd	430	;
		10'd590	:	SINE_TMP	 =	9'd	429	;
		10'd591	:	SINE_TMP	 =	9'd	428	;
		10'd592	:	SINE_TMP	 =	9'd	427	;
		10'd593	:	SINE_TMP	 =	9'd	426	;
		10'd594	:	SINE_TMP	 =	9'd	425	;
		10'd595	:	SINE_TMP	 =	9'd	424	;
		10'd596	:	SINE_TMP	 =	9'd	423	;
		10'd597	:	SINE_TMP	 =	9'd	422	;
		10'd598	:	SINE_TMP	 =	9'd	421	;
		10'd599	:	SINE_TMP	 =	9'd	420	;
		10'd600	:	SINE_TMP	 =	9'd	419	;
		10'd601	:	SINE_TMP	 =	9'd	418	;
		10'd602	:	SINE_TMP	 =	9'd	417	;
		10'd603	:	SINE_TMP	 =	9'd	416	;
		10'd604	:	SINE_TMP	 =	9'd	415	;
		10'd605	:	SINE_TMP	 =	9'd	414	;
		10'd606	:	SINE_TMP	 =	9'd	413	;
		10'd607	:	SINE_TMP	 =	9'd	412	;
		10'd608	:	SINE_TMP	 =	9'd	411	;
		10'd609	:	SINE_TMP	 =	9'd	410	;
		10'd610	:	SINE_TMP	 =	9'd	409	;
		10'd611	:	SINE_TMP	 =	9'd	408	;
		10'd612	:	SINE_TMP	 =	9'd	407	;
		10'd613	:	SINE_TMP	 =	9'd	406	;
		10'd614	:	SINE_TMP	 =	9'd	405	;
		10'd615	:	SINE_TMP	 =	9'd	404	;
		10'd616	:	SINE_TMP	 =	9'd	403	;
		10'd617	:	SINE_TMP	 =	9'd	402	;
		10'd618	:	SINE_TMP	 =	9'd	401	;
		10'd619	:	SINE_TMP	 =	9'd	400	;
		10'd620	:	SINE_TMP	 =	9'd	399	;
		10'd621	:	SINE_TMP	 =	9'd	398	;
		10'd622	:	SINE_TMP	 =	9'd	397	;
		10'd623	:	SINE_TMP	 =	9'd	395	;
		10'd624	:	SINE_TMP	 =	9'd	394	;
		10'd625	:	SINE_TMP	 =	9'd	393	;
		10'd626	:	SINE_TMP	 =	9'd	392	;
		10'd627	:	SINE_TMP	 =	9'd	391	;
		10'd628	:	SINE_TMP	 =	9'd	390	;
		10'd629	:	SINE_TMP	 =	9'd	389	;
		10'd630	:	SINE_TMP	 =	9'd	388	;
		10'd631	:	SINE_TMP	 =	9'd	387	;
		10'd632	:	SINE_TMP	 =	9'd	385	;
		10'd633	:	SINE_TMP	 =	9'd	384	;
		10'd634	:	SINE_TMP	 =	9'd	383	;
		10'd635	:	SINE_TMP	 =	9'd	382	;
		10'd636	:	SINE_TMP	 =	9'd	381	;
		10'd637	:	SINE_TMP	 =	9'd	380	;
		10'd638	:	SINE_TMP	 =	9'd	379	;
		10'd639	:	SINE_TMP	 =	9'd	377	;
		10'd640	:	SINE_TMP	 =	9'd	376	;
		10'd641	:	SINE_TMP	 =	9'd	375	;
		10'd642	:	SINE_TMP	 =	9'd	374	;
		10'd643	:	SINE_TMP	 =	9'd	373	;
		10'd644	:	SINE_TMP	 =	9'd	371	;
		10'd645	:	SINE_TMP	 =	9'd	370	;
		10'd646	:	SINE_TMP	 =	9'd	369	;
		10'd647	:	SINE_TMP	 =	9'd	368	;
		10'd648	:	SINE_TMP	 =	9'd	367	;
		10'd649	:	SINE_TMP	 =	9'd	365	;
		10'd650	:	SINE_TMP	 =	9'd	364	;
		10'd651	:	SINE_TMP	 =	9'd	363	;
		10'd652	:	SINE_TMP	 =	9'd	362	;
		10'd653	:	SINE_TMP	 =	9'd	360	;
		10'd654	:	SINE_TMP	 =	9'd	359	;
		10'd655	:	SINE_TMP	 =	9'd	358	;
		10'd656	:	SINE_TMP	 =	9'd	357	;
		10'd657	:	SINE_TMP	 =	9'd	355	;
		10'd658	:	SINE_TMP	 =	9'd	354	;
		10'd659	:	SINE_TMP	 =	9'd	353	;
		10'd660	:	SINE_TMP	 =	9'd	352	;
		10'd661	:	SINE_TMP	 =	9'd	350	;
		10'd662	:	SINE_TMP	 =	9'd	349	;
		10'd663	:	SINE_TMP	 =	9'd	348	;
		10'd664	:	SINE_TMP	 =	9'd	347	;
		10'd665	:	SINE_TMP	 =	9'd	345	;
		10'd666	:	SINE_TMP	 =	9'd	344	;
		10'd667	:	SINE_TMP	 =	9'd	343	;
		10'd668	:	SINE_TMP	 =	9'd	341	;
		10'd669	:	SINE_TMP	 =	9'd	340	;
		10'd670	:	SINE_TMP	 =	9'd	339	;
		10'd671	:	SINE_TMP	 =	9'd	337	;
		10'd672	:	SINE_TMP	 =	9'd	336	;
		10'd673	:	SINE_TMP	 =	9'd	335	;
		10'd674	:	SINE_TMP	 =	9'd	333	;
		10'd675	:	SINE_TMP	 =	9'd	332	;
		10'd676	:	SINE_TMP	 =	9'd	331	;
		10'd677	:	SINE_TMP	 =	9'd	329	;
		10'd678	:	SINE_TMP	 =	9'd	328	;
		10'd679	:	SINE_TMP	 =	9'd	327	;
		10'd680	:	SINE_TMP	 =	9'd	325	;
		10'd681	:	SINE_TMP	 =	9'd	324	;
		10'd682	:	SINE_TMP	 =	9'd	323	;
		10'd683	:	SINE_TMP	 =	9'd	321	;
		10'd684	:	SINE_TMP	 =	9'd	320	;
		10'd685	:	SINE_TMP	 =	9'd	318	;
		10'd686	:	SINE_TMP	 =	9'd	317	;
		10'd687	:	SINE_TMP	 =	9'd	316	;
		10'd688	:	SINE_TMP	 =	9'd	314	;
		10'd689	:	SINE_TMP	 =	9'd	313	;
		10'd690	:	SINE_TMP	 =	9'd	312	;
		10'd691	:	SINE_TMP	 =	9'd	310	;
		10'd692	:	SINE_TMP	 =	9'd	309	;
		10'd693	:	SINE_TMP	 =	9'd	307	;
		10'd694	:	SINE_TMP	 =	9'd	306	;
		10'd695	:	SINE_TMP	 =	9'd	304	;
		10'd696	:	SINE_TMP	 =	9'd	303	;
		10'd697	:	SINE_TMP	 =	9'd	302	;
		10'd698	:	SINE_TMP	 =	9'd	300	;
		10'd699	:	SINE_TMP	 =	9'd	299	;
		10'd700	:	SINE_TMP	 =	9'd	297	;
		10'd701	:	SINE_TMP	 =	9'd	296	;
		10'd702	:	SINE_TMP	 =	9'd	294	;
		10'd703	:	SINE_TMP	 =	9'd	293	;
		10'd704	:	SINE_TMP	 =	9'd	292	;
		10'd705	:	SINE_TMP	 =	9'd	290	;
		10'd706	:	SINE_TMP	 =	9'd	289	;
		10'd707	:	SINE_TMP	 =	9'd	287	;
		10'd708	:	SINE_TMP	 =	9'd	286	;
		10'd709	:	SINE_TMP	 =	9'd	284	;
		10'd710	:	SINE_TMP	 =	9'd	283	;
		10'd711	:	SINE_TMP	 =	9'd	281	;
		10'd712	:	SINE_TMP	 =	9'd	280	;
		10'd713	:	SINE_TMP	 =	9'd	278	;
		10'd714	:	SINE_TMP	 =	9'd	277	;
		10'd715	:	SINE_TMP	 =	9'd	275	;
		10'd716	:	SINE_TMP	 =	9'd	274	;
		10'd717	:	SINE_TMP	 =	9'd	272	;
		10'd718	:	SINE_TMP	 =	9'd	271	;
		10'd719	:	SINE_TMP	 =	9'd	269	;
		10'd720	:	SINE_TMP	 =	9'd	268	;
		10'd721	:	SINE_TMP	 =	9'd	266	;
		10'd722	:	SINE_TMP	 =	9'd	265	;
		10'd723	:	SINE_TMP	 =	9'd	263	;
		10'd724	:	SINE_TMP	 =	9'd	262	;
		10'd725	:	SINE_TMP	 =	9'd	260	;
		10'd726	:	SINE_TMP	 =	9'd	259	;
		10'd727	:	SINE_TMP	 =	9'd	257	;
		10'd728	:	SINE_TMP	 =	9'd	256	;
		10'd729	:	SINE_TMP	 =	9'd	254	;
		10'd730	:	SINE_TMP	 =	9'd	253	;
		10'd731	:	SINE_TMP	 =	9'd	251	;
		10'd732	:	SINE_TMP	 =	9'd	249	;
		10'd733	:	SINE_TMP	 =	9'd	248	;
		10'd734	:	SINE_TMP	 =	9'd	246	;
		10'd735	:	SINE_TMP	 =	9'd	245	;
		10'd736	:	SINE_TMP	 =	9'd	243	;
		10'd737	:	SINE_TMP	 =	9'd	242	;
		10'd738	:	SINE_TMP	 =	9'd	240	;
		10'd739	:	SINE_TMP	 =	9'd	239	;
		10'd740	:	SINE_TMP	 =	9'd	237	;
		10'd741	:	SINE_TMP	 =	9'd	235	;
		10'd742	:	SINE_TMP	 =	9'd	234	;
		10'd743	:	SINE_TMP	 =	9'd	232	;
		10'd744	:	SINE_TMP	 =	9'd	231	;
		10'd745	:	SINE_TMP	 =	9'd	229	;
		10'd746	:	SINE_TMP	 =	9'd	227	;
		10'd747	:	SINE_TMP	 =	9'd	226	;
		10'd748	:	SINE_TMP	 =	9'd	224	;
		10'd749	:	SINE_TMP	 =	9'd	223	;
		10'd750	:	SINE_TMP	 =	9'd	221	;
		10'd751	:	SINE_TMP	 =	9'd	219	;
		10'd752	:	SINE_TMP	 =	9'd	218	;
		10'd753	:	SINE_TMP	 =	9'd	216	;
		10'd754	:	SINE_TMP	 =	9'd	215	;
		10'd755	:	SINE_TMP	 =	9'd	213	;
		10'd756	:	SINE_TMP	 =	9'd	211	;
		10'd757	:	SINE_TMP	 =	9'd	210	;
		10'd758	:	SINE_TMP	 =	9'd	208	;
		10'd759	:	SINE_TMP	 =	9'd	207	;
		10'd760	:	SINE_TMP	 =	9'd	205	;
		10'd761	:	SINE_TMP	 =	9'd	203	;
		10'd762	:	SINE_TMP	 =	9'd	202	;
		10'd763	:	SINE_TMP	 =	9'd	200	;
		10'd764	:	SINE_TMP	 =	9'd	198	;
		10'd765	:	SINE_TMP	 =	9'd	197	;
		10'd766	:	SINE_TMP	 =	9'd	195	;
		10'd767	:	SINE_TMP	 =	9'd	193	;
		10'd768	:	SINE_TMP	 =	9'd	192	;
		10'd769	:	SINE_TMP	 =	9'd	190	;
		10'd770	:	SINE_TMP	 =	9'd	188	;
		10'd771	:	SINE_TMP	 =	9'd	187	;
		10'd772	:	SINE_TMP	 =	9'd	185	;
		10'd773	:	SINE_TMP	 =	9'd	183	;
		10'd774	:	SINE_TMP	 =	9'd	182	;
		10'd775	:	SINE_TMP	 =	9'd	180	;
		10'd776	:	SINE_TMP	 =	9'd	178	;
		10'd777	:	SINE_TMP	 =	9'd	177	;
		10'd778	:	SINE_TMP	 =	9'd	175	;
		10'd779	:	SINE_TMP	 =	9'd	173	;
		10'd780	:	SINE_TMP	 =	9'd	172	;
		10'd781	:	SINE_TMP	 =	9'd	170	;
		10'd782	:	SINE_TMP	 =	9'd	168	;
		10'd783	:	SINE_TMP	 =	9'd	167	;
		10'd784	:	SINE_TMP	 =	9'd	165	;
		10'd785	:	SINE_TMP	 =	9'd	163	;
		10'd786	:	SINE_TMP	 =	9'd	162	;
		10'd787	:	SINE_TMP	 =	9'd	160	;
		10'd788	:	SINE_TMP	 =	9'd	158	;
		10'd789	:	SINE_TMP	 =	9'd	157	;
		10'd790	:	SINE_TMP	 =	9'd	155	;
		10'd791	:	SINE_TMP	 =	9'd	153	;
		10'd792	:	SINE_TMP	 =	9'd	151	;
		10'd793	:	SINE_TMP	 =	9'd	150	;
		10'd794	:	SINE_TMP	 =	9'd	148	;
		10'd795	:	SINE_TMP	 =	9'd	146	;
		10'd796	:	SINE_TMP	 =	9'd	145	;
		10'd797	:	SINE_TMP	 =	9'd	143	;
		10'd798	:	SINE_TMP	 =	9'd	141	;
		10'd799	:	SINE_TMP	 =	9'd	139	;
		10'd800	:	SINE_TMP	 =	9'd	138	;
		10'd801	:	SINE_TMP	 =	9'd	136	;
		10'd802	:	SINE_TMP	 =	9'd	134	;
		10'd803	:	SINE_TMP	 =	9'd	133	;
		10'd804	:	SINE_TMP	 =	9'd	131	;
		10'd805	:	SINE_TMP	 =	9'd	129	;
		10'd806	:	SINE_TMP	 =	9'd	127	;
		10'd807	:	SINE_TMP	 =	9'd	126	;
		10'd808	:	SINE_TMP	 =	9'd	124	;
		10'd809	:	SINE_TMP	 =	9'd	122	;
		10'd810	:	SINE_TMP	 =	9'd	120	;
		10'd811	:	SINE_TMP	 =	9'd	119	;
		10'd812	:	SINE_TMP	 =	9'd	117	;
		10'd813	:	SINE_TMP	 =	9'd	115	;
		10'd814	:	SINE_TMP	 =	9'd	114	;
		10'd815	:	SINE_TMP	 =	9'd	112	;
		10'd816	:	SINE_TMP	 =	9'd	110	;
		10'd817	:	SINE_TMP	 =	9'd	108	;
		10'd818	:	SINE_TMP	 =	9'd	107	;
		10'd819	:	SINE_TMP	 =	9'd	105	;
		10'd820	:	SINE_TMP	 =	9'd	103	;
		10'd821	:	SINE_TMP	 =	9'd	101	;
		10'd822	:	SINE_TMP	 =	9'd	100	;
		10'd823	:	SINE_TMP	 =	9'd	98	;
		10'd824	:	SINE_TMP	 =	9'd	96	;
		10'd825	:	SINE_TMP	 =	9'd	94	;
		10'd826	:	SINE_TMP	 =	9'd	92	;
		10'd827	:	SINE_TMP	 =	9'd	91	;
		10'd828	:	SINE_TMP	 =	9'd	89	;
		10'd829	:	SINE_TMP	 =	9'd	87	;
		10'd830	:	SINE_TMP	 =	9'd	85	;
		10'd831	:	SINE_TMP	 =	9'd	84	;
		10'd832	:	SINE_TMP	 =	9'd	82	;
		10'd833	:	SINE_TMP	 =	9'd	80	;
		10'd834	:	SINE_TMP	 =	9'd	78	;
		10'd835	:	SINE_TMP	 =	9'd	77	;
		10'd836	:	SINE_TMP	 =	9'd	75	;
		10'd837	:	SINE_TMP	 =	9'd	73	;
		10'd838	:	SINE_TMP	 =	9'd	71	;
		10'd839	:	SINE_TMP	 =	9'd	70	;
		10'd840	:	SINE_TMP	 =	9'd	68	;
		10'd841	:	SINE_TMP	 =	9'd	66	;
		10'd842	:	SINE_TMP	 =	9'd	64	;
		10'd843	:	SINE_TMP	 =	9'd	62	;
		10'd844	:	SINE_TMP	 =	9'd	61	;
		10'd845	:	SINE_TMP	 =	9'd	59	;
		10'd846	:	SINE_TMP	 =	9'd	57	;
		10'd847	:	SINE_TMP	 =	9'd	55	;
		10'd848	:	SINE_TMP	 =	9'd	54	;
		10'd849	:	SINE_TMP	 =	9'd	52	;
		10'd850	:	SINE_TMP	 =	9'd	50	;
		10'd851	:	SINE_TMP	 =	9'd	48	;
		10'd852	:	SINE_TMP	 =	9'd	46	;
		10'd853	:	SINE_TMP	 =	9'd	45	;
		10'd854	:	SINE_TMP	 =	9'd	43	;
		10'd855	:	SINE_TMP	 =	9'd	41	;
		10'd856	:	SINE_TMP	 =	9'd	39	;
		10'd857	:	SINE_TMP	 =	9'd	38	;
		10'd858	:	SINE_TMP	 =	9'd	36	;
		10'd859	:	SINE_TMP	 =	9'd	34	;
		10'd860	:	SINE_TMP	 =	9'd	32	;
		10'd861	:	SINE_TMP	 =	9'd	30	;
		10'd862	:	SINE_TMP	 =	9'd	29	;
		10'd863	:	SINE_TMP	 =	9'd	27	;
		10'd864	:	SINE_TMP	 =	9'd	25	;
		10'd865	:	SINE_TMP	 =	9'd	23	;
		10'd866	:	SINE_TMP	 =	9'd	21	;
		10'd867	:	SINE_TMP	 =	9'd	20	;
		10'd868	:	SINE_TMP	 =	9'd	18	;
		10'd869	:	SINE_TMP	 =	9'd	16	;
		10'd870	:	SINE_TMP	 =	9'd	14	;
		10'd871	:	SINE_TMP	 =	9'd	13	;
		10'd872	:	SINE_TMP	 =	9'd	11	;
		10'd873	:	SINE_TMP	 =	9'd	9	;
		10'd874	:	SINE_TMP	 =	9'd	7	;
		10'd875	:	SINE_TMP	 =	9'd	5	;
		10'd876	:	SINE_TMP	 =	9'd	4	;
		10'd877	:	SINE_TMP	 =	9'd	2	;
		10'd878	:	SINE_TMP	 =	9'd	0	;
		default: SINE_TMP = 9'd0;
		
	endcase
	SINE_OUT = SINE_TMP;
end
	 

endmodule
