module  sine_look_up(
		input  [8:0] teth_ta,
		//input  clk,
		output reg [10:0] sine_out);
		 
always @(teth_ta) begin      // sine look up table 
	case (teth_ta)                    			
		9'd0	:	sine_out	 =	11'd	0	;
		9'd1	:	sine_out	 =	11'd	24	;
		9'd2	:	sine_out	 =	11'd	48	;
		9'd3	:	sine_out	 =	11'd	72	;
		9'd4	:	sine_out	 =	11'd	95	;
		9'd5	:	sine_out	 =	11'd	119	;
		9'd6	:	sine_out	 =	11'd	143	;
		9'd7	:	sine_out	 =	11'd	167	;
		9'd8	:	sine_out	 =	11'd	191	;
		9'd9	:	sine_out	 =	11'd	214	;
		9'd10	:	sine_out	 =	11'd	238	;
		9'd11	:	sine_out	 =	11'd	262	;
		9'd12	:	sine_out	 =	11'd	285	;
		9'd13	:	sine_out	 =	11'd	309	;
		9'd14	:	sine_out	 =	11'd	333	;
		9'd15	:	sine_out	 =	11'd	356	;
		9'd16	:	sine_out	 =	11'd	379	;
		9'd17	:	sine_out	 =	11'd	403	;
		9'd18	:	sine_out	 =	11'd	426	;
		9'd19	:	sine_out	 =	11'd	449	;
		9'd20	:	sine_out	 =	11'd	473	;
		9'd21	:	sine_out	 =	11'd	496	;
		9'd22	:	sine_out	 =	11'd	519	;
		9'd23	:	sine_out	 =	11'd	542	;
		9'd24	:	sine_out	 =	11'd	564	;
		9'd25	:	sine_out	 =	11'd	587	;
		9'd26	:	sine_out	 =	11'd	610	;
		9'd27	:	sine_out	 =	11'd	632	;
		9'd28	:	sine_out	 =	11'd	655	;
		9'd29	:	sine_out	 =	11'd	677	;
		9'd30	:	sine_out	 =	11'd	699	;
		9'd31	:	sine_out	 =	11'd	722	;
		9'd32	:	sine_out	 =	11'd	744	;
		9'd33	:	sine_out	 =	11'd	766	;
		9'd34	:	sine_out	 =	11'd	787	;
		9'd35	:	sine_out	 =	11'd	809	;
		9'd36	:	sine_out	 =	11'd	831	;
		9'd37	:	sine_out	 =	11'd	852	;
		9'd38	:	sine_out	 =	11'd	873	;
		9'd39	:	sine_out	 =	11'd	894	;
		9'd40	:	sine_out	 =	11'd	915	;
		9'd41	:	sine_out	 =	11'd	936	;
		9'd42	:	sine_out	 =	11'd	957	;
		9'd43	:	sine_out	 =	11'd	977	;
		9'd44	:	sine_out	 =	11'd	998	;
		9'd45	:	sine_out	 =	11'd	1018	;
		9'd46	:	sine_out	 =	11'd	1038	;
		9'd47	:	sine_out	 =	11'd	1058	;
		9'd48	:	sine_out	 =	11'd	1078	;
		9'd49	:	sine_out	 =	11'd	1097	;
		9'd50	:	sine_out	 =	11'd	1117	;
		9'd51	:	sine_out	 =	11'd	1136	;
		9'd52	:	sine_out	 =	11'd	1155	;
		9'd53	:	sine_out	 =	11'd	1174	;
		9'd54	:	sine_out	 =	11'd	1193	;
		9'd55	:	sine_out	 =	11'd	1211	;
		9'd56	:	sine_out	 =	11'd	1229	;
		9'd57	:	sine_out	 =	11'd	1248	;
		9'd58	:	sine_out	 =	11'd	1265	;
		9'd59	:	sine_out	 =	11'd	1283	;
		9'd60	:	sine_out	 =	11'd	1301	;
		9'd61	:	sine_out	 =	11'd	1318	;
		9'd62	:	sine_out	 =	11'd	1335	;
		9'd63	:	sine_out	 =	11'd	1352	;
		9'd64	:	sine_out	 =	11'd	1369	;
		9'd65	:	sine_out	 =	11'd	1385	;
		9'd66	:	sine_out	 =	11'd	1401	;
		9'd67	:	sine_out	 =	11'd	1417	;
		9'd68	:	sine_out	 =	11'd	1433	;
		9'd69	:	sine_out	 =	11'd	1449	;
		9'd70	:	sine_out	 =	11'd	1464	;
		9'd71	:	sine_out	 =	11'd	1479	;
		9'd72	:	sine_out	 =	11'd	1494	;
		9'd73	:	sine_out	 =	11'd	1509	;
		9'd74	:	sine_out	 =	11'd	1523	;
		9'd75	:	sine_out	 =	11'd	1537	;
		9'd76	:	sine_out	 =	11'd	1551	;
		9'd77	:	sine_out	 =	11'd	1565	;
		9'd78	:	sine_out	 =	11'd	1578	;
		9'd79	:	sine_out	 =	11'd	1591	;
		9'd80	:	sine_out	 =	11'd	1604	;
		9'd81	:	sine_out	 =	11'd	1617	;
		9'd82	:	sine_out	 =	11'd	1629	;
		9'd83	:	sine_out	 =	11'd	1641	;
		9'd84	:	sine_out	 =	11'd	1653	;
		9'd85	:	sine_out	 =	11'd	1665	;
		9'd86	:	sine_out	 =	11'd	1676	;
		9'd87	:	sine_out	 =	11'd	1687	;
		9'd88	:	sine_out	 =	11'd	1698	;
		9'd89	:	sine_out	 =	11'd	1709	;
		9'd90	:	sine_out	 =	11'd	1719	;
		9'd91	:	sine_out	 =	11'd	1729	;
		9'd92	:	sine_out	 =	11'd	1739	;
		9'd93	:	sine_out	 =	11'd	1748	;
		9'd94	:	sine_out	 =	11'd	1758	;
		9'd95	:	sine_out	 =	11'd	1767	;
		9'd96	:	sine_out	 =	11'd	1775	;
		9'd97	:	sine_out	 =	11'd	1784	;
		9'd98	:	sine_out	 =	11'd	1792	;
		9'd99	:	sine_out	 =	11'd	1799	;
		9'd100	:	sine_out	 =	11'd	1807	;
		9'd101	:	sine_out	 =	11'd	1814	;
		9'd102	:	sine_out	 =	11'd	1821	;
		9'd103	:	sine_out	 =	11'd	1828	;
		9'd104	:	sine_out	 =	11'd	1834	;
		9'd105	:	sine_out	 =	11'd	1840	;
		9'd106	:	sine_out	 =	11'd	1846	;
		9'd107	:	sine_out	 =	11'd	1852	;
		9'd108	:	sine_out	 =	11'd	1857	;
		9'd109	:	sine_out	 =	11'd	1862	;
		9'd110	:	sine_out	 =	11'd	1866	;
		9'd111	:	sine_out	 =	11'd	1871	;
		9'd112	:	sine_out	 =	11'd	1875	;
		9'd113	:	sine_out	 =	11'd	1878	;
		9'd114	:	sine_out	 =	11'd	1882	;
		9'd115	:	sine_out	 =	11'd	1885	;
		9'd116	:	sine_out	 =	11'd	1888	;
		9'd117	:	sine_out	 =	11'd	1890	;
		9'd118	:	sine_out	 =	11'd	1893	;
		9'd119	:	sine_out	 =	11'd	1895	;
		9'd120	:	sine_out	 =	11'd	1896	;
		9'd121	:	sine_out	 =	11'd	1898	;
		9'd122	:	sine_out	 =	11'd	1899	;
		9'd123	:	sine_out	 =	11'd	1899	;
		9'd124	:	sine_out	 =	11'd	1900	;
		9'd125	:	sine_out	 =	11'd	1900	;
		9'd126	:	sine_out	 =	11'd	1900	;
		9'd127	:	sine_out	 =	11'd	1899	;
		9'd128	:	sine_out	 =	11'd	1899	;
		9'd129	:	sine_out	 =	11'd	1898	;
		9'd130	:	sine_out	 =	11'd	1896	;
		9'd131	:	sine_out	 =	11'd	1895	;
		9'd132	:	sine_out	 =	11'd	1893	;
		9'd133	:	sine_out	 =	11'd	1890	;
		9'd134	:	sine_out	 =	11'd	1888	;
		9'd135	:	sine_out	 =	11'd	1885	;
		9'd136	:	sine_out	 =	11'd	1882	;
		9'd137	:	sine_out	 =	11'd	1878	;
		9'd138	:	sine_out	 =	11'd	1875	;
		9'd139	:	sine_out	 =	11'd	1871	;
		9'd140	:	sine_out	 =	11'd	1866	;
		9'd141	:	sine_out	 =	11'd	1862	;
		9'd142	:	sine_out	 =	11'd	1857	;
		9'd143	:	sine_out	 =	11'd	1852	;
		9'd144	:	sine_out	 =	11'd	1846	;
		9'd145	:	sine_out	 =	11'd	1840	;
		9'd146	:	sine_out	 =	11'd	1834	;
		9'd147	:	sine_out	 =	11'd	1828	;
		9'd148	:	sine_out	 =	11'd	1821	;
		9'd149	:	sine_out	 =	11'd	1814	;
		9'd150	:	sine_out	 =	11'd	1807	;
		9'd151	:	sine_out	 =	11'd	1799	;
		9'd152	:	sine_out	 =	11'd	1792	;
		9'd153	:	sine_out	 =	11'd	1784	;
		9'd154	:	sine_out	 =	11'd	1775	;
		9'd155	:	sine_out	 =	11'd	1767	;
		9'd156	:	sine_out	 =	11'd	1758	;
		9'd157	:	sine_out	 =	11'd	1748	;
		9'd158	:	sine_out	 =	11'd	1739	;
		9'd159	:	sine_out	 =	11'd	1729	;
		9'd160	:	sine_out	 =	11'd	1719	;
		9'd161	:	sine_out	 =	11'd	1709	;
		9'd162	:	sine_out	 =	11'd	1698	;
		9'd163	:	sine_out	 =	11'd	1687	;
		9'd164	:	sine_out	 =	11'd	1676	;
		9'd165	:	sine_out	 =	11'd	1665	;
		9'd166	:	sine_out	 =	11'd	1653	;
		9'd167	:	sine_out	 =	11'd	1641	;
		9'd168	:	sine_out	 =	11'd	1629	;
		9'd169	:	sine_out	 =	11'd	1617	;
		9'd170	:	sine_out	 =	11'd	1604	;
		9'd171	:	sine_out	 =	11'd	1591	;
		9'd172	:	sine_out	 =	11'd	1578	;
		9'd173	:	sine_out	 =	11'd	1565	;
		9'd174	:	sine_out	 =	11'd	1551	;
		9'd175	:	sine_out	 =	11'd	1537	;
		9'd176	:	sine_out	 =	11'd	1523	;
		9'd177	:	sine_out	 =	11'd	1509	;
		9'd178	:	sine_out	 =	11'd	1494	;
		9'd179	:	sine_out	 =	11'd	1479	;
		9'd180	:	sine_out	 =	11'd	1464	;
		9'd181	:	sine_out	 =	11'd	1449	;
		9'd182	:	sine_out	 =	11'd	1433	;
		9'd183	:	sine_out	 =	11'd	1417	;
		9'd184	:	sine_out	 =	11'd	1401	;
		9'd185	:	sine_out	 =	11'd	1385	;
		9'd186	:	sine_out	 =	11'd	1369	;
		9'd187	:	sine_out	 =	11'd	1352	;
		9'd188	:	sine_out	 =	11'd	1335	;
		9'd189	:	sine_out	 =	11'd	1318	;
		9'd190	:	sine_out	 =	11'd	1301	;
		9'd191	:	sine_out	 =	11'd	1283	;
		9'd192	:	sine_out	 =	11'd	1265	;
		9'd193	:	sine_out	 =	11'd	1248	;
		9'd194	:	sine_out	 =	11'd	1229	;
		9'd195	:	sine_out	 =	11'd	1211	;
		9'd196	:	sine_out	 =	11'd	1193	;
		9'd197	:	sine_out	 =	11'd	1174	;
		9'd198	:	sine_out	 =	11'd	1155	;
		9'd199	:	sine_out	 =	11'd	1136	;
		9'd200	:	sine_out	 =	11'd	1117	;
		9'd201	:	sine_out	 =	11'd	1097	;
		9'd202	:	sine_out	 =	11'd	1078	;
		9'd203	:	sine_out	 =	11'd	1058	;
		9'd204	:	sine_out	 =	11'd	1038	;
		9'd205	:	sine_out	 =	11'd	1018	;
		9'd206	:	sine_out	 =	11'd	998	;
		9'd207	:	sine_out	 =	11'd	977	;
		9'd208	:	sine_out	 =	11'd	957	;
		9'd209	:	sine_out	 =	11'd	936	;
		9'd210	:	sine_out	 =	11'd	915	;
		9'd211	:	sine_out	 =	11'd	894	;
		9'd212	:	sine_out	 =	11'd	873	;
		9'd213	:	sine_out	 =	11'd	852	;
		9'd214	:	sine_out	 =	11'd	831	;
		9'd215	:	sine_out	 =	11'd	809	;
		9'd216	:	sine_out	 =	11'd	787	;
		9'd217	:	sine_out	 =	11'd	766	;
		9'd218	:	sine_out	 =	11'd	744	;
		9'd219	:	sine_out	 =	11'd	722	;
		9'd220	:	sine_out	 =	11'd	699	;
		9'd221	:	sine_out	 =	11'd	677	;
		9'd222	:	sine_out	 =	11'd	655	;
		9'd223	:	sine_out	 =	11'd	632	;
		9'd224	:	sine_out	 =	11'd	610	;
		9'd225	:	sine_out	 =	11'd	587	;
		9'd226	:	sine_out	 =	11'd	564	;
		9'd227	:	sine_out	 =	11'd	542	;
		9'd228	:	sine_out	 =	11'd	519	;
		9'd229	:	sine_out	 =	11'd	496	;
		9'd230	:	sine_out	 =	11'd	473	;
		9'd231	:	sine_out	 =	11'd	449	;
		9'd232	:	sine_out	 =	11'd	426	;
		9'd233	:	sine_out	 =	11'd	403	;
		9'd234	:	sine_out	 =	11'd	379	;
		9'd235	:	sine_out	 =	11'd	356	;
		9'd236	:	sine_out	 =	11'd	333	;
		9'd237	:	sine_out	 =	11'd	309	;
		9'd238	:	sine_out	 =	11'd	285	;
		9'd239	:	sine_out	 =	11'd	262	;
		9'd240	:	sine_out	 =	11'd	238	;
		9'd241	:	sine_out	 =	11'd	214	;
		9'd242	:	sine_out	 =	11'd	191	;
		9'd243	:	sine_out	 =	11'd	167	;
		9'd244	:	sine_out	 =	11'd	143	;
		9'd245	:	sine_out	 =	11'd	119	;
		9'd246	:	sine_out	 =	11'd	95	;
		9'd247	:	sine_out	 =	11'd	72	;
		9'd248	:	sine_out	 =	11'd	48	;
		9'd249	:	sine_out	 =	11'd	24	;
		9'd250	:	sine_out	 =	11'd	0	;
		9'd251	:	sine_out	 =	11'd	0	;
		9'd252	:	sine_out	 =	11'd	0	;
		9'd253	:	sine_out	 =	11'd	0	;
		9'd254	:	sine_out	 =	11'd	0	;
		9'd255	:	sine_out	 =	11'd	0	;
		9'd256	:	sine_out	 =	11'd	0	;
		9'd257	:	sine_out	 =	11'd	0	;
		9'd258	:	sine_out	 =	11'd	0	;
		9'd259	:	sine_out	 =	11'd	0	;
		9'd260	:	sine_out	 =	11'd	0	;
		9'd261	:	sine_out	 =	11'd	0	;
		9'd262	:	sine_out	 =	11'd	0	;
		9'd263	:	sine_out	 =	11'd	0	;
		9'd264	:	sine_out	 =	11'd	0	;
		9'd265	:	sine_out	 =	11'd	0	;
		9'd266	:	sine_out	 =	11'd	0	;
		9'd267	:	sine_out	 =	11'd	0	;
		9'd268	:	sine_out	 =	11'd	0	;
		9'd269	:	sine_out	 =	11'd	0	;
		9'd270	:	sine_out	 =	11'd	0	;
		9'd271	:	sine_out	 =	11'd	0	;
		9'd272	:	sine_out	 =	11'd	0	;
		9'd273	:	sine_out	 =	11'd	0	;
		9'd274	:	sine_out	 =	11'd	0	;
		9'd275	:	sine_out	 =	11'd	0	;
		9'd276	:	sine_out	 =	11'd	0	;
		9'd277	:	sine_out	 =	11'd	0	;
		9'd278	:	sine_out	 =	11'd	0	;
		9'd279	:	sine_out	 =	11'd	0	;
		9'd280	:	sine_out	 =	11'd	0	;
		9'd281	:	sine_out	 =	11'd	0	;
		9'd282	:	sine_out	 =	11'd	0	;
		9'd283	:	sine_out	 =	11'd	0	;
		9'd284	:	sine_out	 =	11'd	0	;
		9'd285	:	sine_out	 =	11'd	0	;
		9'd286	:	sine_out	 =	11'd	0	;
		9'd287	:	sine_out	 =	11'd	0	;
		9'd288	:	sine_out	 =	11'd	0	;
		9'd289	:	sine_out	 =	11'd	0	;
		9'd290	:	sine_out	 =	11'd	0	;
		9'd291	:	sine_out	 =	11'd	0	;
		9'd292	:	sine_out	 =	11'd	0	;
		9'd293	:	sine_out	 =	11'd	0	;
		9'd294	:	sine_out	 =	11'd	0	;
		9'd295	:	sine_out	 =	11'd	0	;
		9'd296	:	sine_out	 =	11'd	0	;
		9'd297	:	sine_out	 =	11'd	0	;
		9'd298	:	sine_out	 =	11'd	0	;
		9'd299	:	sine_out	 =	11'd	0	;
		9'd300	:	sine_out	 =	11'd	0	;
		9'd301	:	sine_out	 =	11'd	0	;
		9'd302	:	sine_out	 =	11'd	0	;
		9'd303	:	sine_out	 =	11'd	0	;
		9'd304	:	sine_out	 =	11'd	0	;
		9'd305	:	sine_out	 =	11'd	0	;
		9'd306	:	sine_out	 =	11'd	0	;
		9'd307	:	sine_out	 =	11'd	0	;
		9'd308	:	sine_out	 =	11'd	0	;
		9'd309	:	sine_out	 =	11'd	0	;
		9'd310	:	sine_out	 =	11'd	0	;
		9'd311	:	sine_out	 =	11'd	0	;
		9'd312	:	sine_out	 =	11'd	0	;
		9'd313	:	sine_out	 =	11'd	0	;
		9'd314	:	sine_out	 =	11'd	0	;
		9'd315	:	sine_out	 =	11'd	0	;
		9'd316	:	sine_out	 =	11'd	0	;
		9'd317	:	sine_out	 =	11'd	0	;
		9'd318	:	sine_out	 =	11'd	0	;
		9'd319	:	sine_out	 =	11'd	0	;
		9'd320	:	sine_out	 =	11'd	0	;
		9'd321	:	sine_out	 =	11'd	0	;
		9'd322	:	sine_out	 =	11'd	0	;
		9'd323	:	sine_out	 =	11'd	0	;
		9'd324	:	sine_out	 =	11'd	0	;
		9'd325	:	sine_out	 =	11'd	0	;
		9'd326	:	sine_out	 =	11'd	0	;
		9'd327	:	sine_out	 =	11'd	0	;
		9'd328	:	sine_out	 =	11'd	0	;
		9'd329	:	sine_out	 =	11'd	0	;
		9'd330	:	sine_out	 =	11'd	0	;
		9'd331	:	sine_out	 =	11'd	0	;
		9'd332	:	sine_out	 =	11'd	0	;
		9'd333	:	sine_out	 =	11'd	0	;
		9'd334	:	sine_out	 =	11'd	0	;
		9'd335	:	sine_out	 =	11'd	0	;
		9'd336	:	sine_out	 =	11'd	0	;
		9'd337	:	sine_out	 =	11'd	0	;
		9'd338	:	sine_out	 =	11'd	0	;
		9'd339	:	sine_out	 =	11'd	0	;
		9'd340	:	sine_out	 =	11'd	0	;
		9'd341	:	sine_out	 =	11'd	0	;
		9'd342	:	sine_out	 =	11'd	0	;
		9'd343	:	sine_out	 =	11'd	0	;
		9'd344	:	sine_out	 =	11'd	0	;
		9'd345	:	sine_out	 =	11'd	0	;
		9'd346	:	sine_out	 =	11'd	0	;
		9'd347	:	sine_out	 =	11'd	0	;
		9'd348	:	sine_out	 =	11'd	0	;
		9'd349	:	sine_out	 =	11'd	0	;
		9'd350	:	sine_out	 =	11'd	0	;
		9'd351	:	sine_out	 =	11'd	0	;
		9'd352	:	sine_out	 =	11'd	0	;
		9'd353	:	sine_out	 =	11'd	0	;
		9'd354	:	sine_out	 =	11'd	0	;
		9'd355	:	sine_out	 =	11'd	0	;
		9'd356	:	sine_out	 =	11'd	0	;
		9'd357	:	sine_out	 =	11'd	0	;
		9'd358	:	sine_out	 =	11'd	0	;
		9'd359	:	sine_out	 =	11'd	0	;
		9'd360	:	sine_out	 =	11'd	0	;
		9'd361	:	sine_out	 =	11'd	0	;
		9'd362	:	sine_out	 =	11'd	0	;
		9'd363	:	sine_out	 =	11'd	0	;
		9'd364	:	sine_out	 =	11'd	0	;
		9'd365	:	sine_out	 =	11'd	0	;
		9'd366	:	sine_out	 =	11'd	0	;
		9'd367	:	sine_out	 =	11'd	0	;
		9'd368	:	sine_out	 =	11'd	0	;
		9'd369	:	sine_out	 =	11'd	0	;
		9'd370	:	sine_out	 =	11'd	0	;
		9'd371	:	sine_out	 =	11'd	0	;
		9'd372	:	sine_out	 =	11'd	0	;
		9'd373	:	sine_out	 =	11'd	0	;
		9'd374	:	sine_out	 =	11'd	0	;
		9'd375	:	sine_out	 =	11'd	0	;
		9'd376	:	sine_out	 =	11'd	0	;
		9'd377	:	sine_out	 =	11'd	0	;
		9'd378	:	sine_out	 =	11'd	0	;
		9'd379	:	sine_out	 =	11'd	0	;
		9'd380	:	sine_out	 =	11'd	0	;
		9'd381	:	sine_out	 =	11'd	0	;
		9'd382	:	sine_out	 =	11'd	0	;
		9'd383	:	sine_out	 =	11'd	0	;
		9'd384	:	sine_out	 =	11'd	0	;
		9'd385	:	sine_out	 =	11'd	0	;
		9'd386	:	sine_out	 =	11'd	0	;
		9'd387	:	sine_out	 =	11'd	0	;
		9'd388	:	sine_out	 =	11'd	0	;
		9'd389	:	sine_out	 =	11'd	0	;
		9'd390	:	sine_out	 =	11'd	0	;
		9'd391	:	sine_out	 =	11'd	0	;
		9'd392	:	sine_out	 =	11'd	0	;
		9'd393	:	sine_out	 =	11'd	0	;
		9'd394	:	sine_out	 =	11'd	0	;
		9'd395	:	sine_out	 =	11'd	0	;
		9'd396	:	sine_out	 =	11'd	0	;
		9'd397	:	sine_out	 =	11'd	0	;
		9'd398	:	sine_out	 =	11'd	0	;
		9'd399	:	sine_out	 =	11'd	0	;
		9'd400	:	sine_out	 =	11'd	0	;
		9'd401	:	sine_out	 =	11'd	0	;
		9'd402	:	sine_out	 =	11'd	0	;
		9'd403	:	sine_out	 =	11'd	0	;
		9'd404	:	sine_out	 =	11'd	0	;
		9'd405	:	sine_out	 =	11'd	0	;
		9'd406	:	sine_out	 =	11'd	0	;
		9'd407	:	sine_out	 =	11'd	0	;
		9'd408	:	sine_out	 =	11'd	0	;
		9'd409	:	sine_out	 =	11'd	0	;
		9'd410	:	sine_out	 =	11'd	0	;
		9'd411	:	sine_out	 =	11'd	0	;
		9'd412	:	sine_out	 =	11'd	0	;
		9'd413	:	sine_out	 =	11'd	0	;
		9'd414	:	sine_out	 =	11'd	0	;
		9'd415	:	sine_out	 =	11'd	0	;
		9'd416	:	sine_out	 =	11'd	0	;
		9'd417	:	sine_out	 =	11'd	0	;
		9'd418	:	sine_out	 =	11'd	0	;
		9'd419	:	sine_out	 =	11'd	0	;
		9'd420	:	sine_out	 =	11'd	0	;
		9'd421	:	sine_out	 =	11'd	0	;
		9'd422	:	sine_out	 =	11'd	0	;
		9'd423	:	sine_out	 =	11'd	0	;
		9'd424	:	sine_out	 =	11'd	0	;
		9'd425	:	sine_out	 =	11'd	0	;
		9'd426	:	sine_out	 =	11'd	0	;
		9'd427	:	sine_out	 =	11'd	0	;
		9'd428	:	sine_out	 =	11'd	0	;
		9'd429	:	sine_out	 =	11'd	0	;
		9'd430	:	sine_out	 =	11'd	0	;
		9'd431	:	sine_out	 =	11'd	0	;
		9'd432	:	sine_out	 =	11'd	0	;
		9'd433	:	sine_out	 =	11'd	0	;
		9'd434	:	sine_out	 =	11'd	0	;
		9'd435	:	sine_out	 =	11'd	0	;
		9'd436	:	sine_out	 =	11'd	0	;
		9'd437	:	sine_out	 =	11'd	0	;
		9'd438	:	sine_out	 =	11'd	0	;
		9'd439	:	sine_out	 =	11'd	0	;
		9'd440	:	sine_out	 =	11'd	0	;
		9'd441	:	sine_out	 =	11'd	0	;
		9'd442	:	sine_out	 =	11'd	0	;
		9'd443	:	sine_out	 =	11'd	0	;
		9'd444	:	sine_out	 =	11'd	0	;
		9'd445	:	sine_out	 =	11'd	0	;
		9'd446	:	sine_out	 =	11'd	0	;
		9'd447	:	sine_out	 =	11'd	0	;
		9'd448	:	sine_out	 =	11'd	0	;
		9'd449	:	sine_out	 =	11'd	0	;
		9'd450	:	sine_out	 =	11'd	0	;
		9'd451	:	sine_out	 =	11'd	0	;
		9'd452	:	sine_out	 =	11'd	0	;
		9'd453	:	sine_out	 =	11'd	0	;
		9'd454	:	sine_out	 =	11'd	0	;
		9'd455	:	sine_out	 =	11'd	0	;
		9'd456	:	sine_out	 =	11'd	0	;
		9'd457	:	sine_out	 =	11'd	0	;
		9'd458	:	sine_out	 =	11'd	0	;
		9'd459	:	sine_out	 =	11'd	0	;
		9'd460	:	sine_out	 =	11'd	0	;
		9'd461	:	sine_out	 =	11'd	0	;
		9'd462	:	sine_out	 =	11'd	0	;
		9'd463	:	sine_out	 =	11'd	0	;
		9'd464	:	sine_out	 =	11'd	0	;
		9'd465	:	sine_out	 =	11'd	0	;
		9'd466	:	sine_out	 =	11'd	0	;
		9'd467	:	sine_out	 =	11'd	0	;
		9'd468	:	sine_out	 =	11'd	0	;
		9'd469	:	sine_out	 =	11'd	0	;
		9'd470	:	sine_out	 =	11'd	0	;
		9'd471	:	sine_out	 =	11'd	0	;
		9'd472	:	sine_out	 =	11'd	0	;
		9'd473	:	sine_out	 =	11'd	0	;
		9'd474	:	sine_out	 =	11'd	0	;
		9'd475	:	sine_out	 =	11'd	0	;
		9'd476	:	sine_out	 =	11'd	0	;
		9'd477	:	sine_out	 =	11'd	0	;
		9'd478	:	sine_out	 =	11'd	0	;
		9'd479	:	sine_out	 =	11'd	0	;
		9'd480	:	sine_out	 =	11'd	0	;
		9'd481	:	sine_out	 =	11'd	0	;
		9'd482	:	sine_out	 =	11'd	0	;
		9'd483	:	sine_out	 =	11'd	0	;
		9'd484	:	sine_out	 =	11'd	0	;
		9'd485	:	sine_out	 =	11'd	0	;
		9'd486	:	sine_out	 =	11'd	0	;
		9'd487	:	sine_out	 =	11'd	0	;
		9'd488	:	sine_out	 =	11'd	0	;
		9'd489	:	sine_out	 =	11'd	0	;
		9'd490	:	sine_out	 =	11'd	0	;
		9'd491	:	sine_out	 =	11'd	0	;
		9'd492	:	sine_out	 =	11'd	0	;
		9'd493	:	sine_out	 =	11'd	0	;
		9'd494	:	sine_out	 =	11'd	0	;
		9'd495	:	sine_out	 =	11'd	0	;
		9'd496	:	sine_out	 =	11'd	0	;
		9'd497	:	sine_out	 =	11'd	0	;
		9'd498	:	sine_out	 =	11'd	0	;
		9'd499	:	sine_out	 =	11'd	0	;



		default: sine_out = 11'd0;
		
	endcase
	
end
endmodule
